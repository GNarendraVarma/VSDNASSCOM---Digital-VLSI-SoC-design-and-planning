* SPICE3 file created from sky130_inv.ext - technology: sky130A

.option scale=0.01u
.include ./libs/pshort.lib
.include ./libs/nshort.lib

//.subckt sky130_inv A Y VPWR VGND
M1000 Y A VPWR VPWR pshort_model.0 w=37 l=23
+ ad=1443 pd=152 as=1517 ps=156
M1001 Y A VGND VGND nshort_model.0 w=35 l=23
+ ad=1435 pd=152 as=1365 ps=148

VDD VPWR 0 3.3V
VSS VGND 0 0V

Va A VGND PULSE(0V 3.3V 0 0.1ns 0.1ns 2ns 4ns)
C0 A Y 0.85f
C1 Y VPWR 0.11f
C2 Y VPWR 0.07f
C3 Y 0 2f
C4 VPWR 0 0.59f
//.ends

.tran 1n 20n
.control
run
.endc
.end


